CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 71 960 1050
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
93 D:\university\semestr.03\Electronics\_���������_�����������\CM60_RUS_ENG\CM60_RUS_ENG\BOM.DAT
0 7
0 71 960 1050
144179219 0
0
6 Title:
5 Name:
0
0
0
6
7 Ground~
168 398 441 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
11 Signal Gen~
195 281 340 0 19 64
0 4 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1065353216
20
1 1000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -1/1V
-18 -30 17 -22
2 V1
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(0 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
4441 0 0
0
0
10 Capacitor~
219 434 318 0 2 5
0 5 3
0
0 0 848 0
3 5uF
-11 -18 10 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3618 0 0
0
0
9 Inductor~
219 408 271 0 2 5
0 4 3
0
0 0 848 0
3 6mH
-11 -17 10 -9
2 L1
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
6153 0 0
0
0
11 Resistor:A~
219 478 358 0 3 5
0 2 3 -1
0
0 0 880 90
1 5
11 0 18 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5394 0 0
0
0
11 Resistor:A~
219 376 318 0 2 5
0 4 5
0
0 0 880 0
2 10
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7734 0 0
0
0
7
2 0 3 0 0 8320 0 4 0 0 6 3
426 271
461 271
461 318
1 0 4 0 0 4224 0 4 0 0 5 3
390 271
338 271
338 318
1 0 2 0 0 4096 0 1 0 0 4 2
398 435
398 386
2 1 2 0 0 12416 0 2 5 0 0 5
312 345
319 345
319 386
478 386
478 376
1 1 4 0 0 0 0 2 6 0 0 4
312 335
320 335
320 318
358 318
2 2 3 0 0 0 0 3 5 0 0 3
443 318
478 318
478 340
2 1 5 0 0 4224 0 6 3 0 0 2
394 318
425 318
0
0
24 0 1
0
0
0
0 0 0
0
0 0 0
1000 0 1 50000
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
1182144 8550464 100 100 0 0
77 66 917 396
960 71 1920 560
917 66
77 66
917 66
917 396
0 0
0.005 0 1.2 -1.2 0.005 0.005
12401 0
4 0.001 0.5
2
331 318
0 4 0 0 3	0 5 0 0
478 321
0 3 0 0 2	0 6 0 0
1051000 4356170 100 100 0 0
77 66 917 396
960 560 1920 1049
568 66
77 66
927 66
927 341
0 0
774.794 1 0.8 -1.2 49999 49999
12387 0
4 1 2
2
327 318
0 4 0 0 3	0 5 0 0
478 325
0 3 0 0 2	0 6 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
