CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 71 960 1050
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
107 Z:\mnt\sda3\Downloads\Firefox\���������_�����������\���������_�����������\CM60_RUS_ENG\CM60_RUS_ENG\BOM.DAT
0 7
0 71 960 1050
144179219 0
0
6 Title:
5 Name:
0
0
0
6
11 Signal Gen~
195 424 285 0 19 64
0 4 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1065353216
20
1 1000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -1/1V
-18 -30 17 -22
2 V1
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(0 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
8953 0 0
0
0
7 Ground~
168 573 346 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4441 0 0
0
0
10 Capacitor~
219 642 285 0 2 5
0 2 3
0
0 0 848 90
5 6.8nF
4 0 39 8
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3618 0 0
0
0
10 Capacitor~
219 525 251 0 2 5
0 4 5
0
0 0 848 0
4 10nF
-14 -18 14 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6153 0 0
0
0
11 Resistor:A~
219 693 286 0 3 5
0 2 3 -1
0
0 0 880 90
2 1G
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5394 0 0
0
0
11 Resistor:A~
219 589 251 0 2 5
0 5 3
0
0 0 880 0
4 100k
-14 -14 14 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7734 0 0
0
0
7
1 0 2 0 0 8192 0 5 0 0 5 3
693 304
693 310
642 310
0 2 3 0 0 4224 0 0 5 6 0 3
642 251
693 251
693 268
1 0 2 0 0 0 0 2 0 0 5 2
573 340
573 311
1 1 4 0 0 4224 0 4 1 0 0 4
516 251
463 251
463 280
455 280
1 2 2 0 0 8320 0 3 1 0 0 5
642 294
642 311
463 311
463 290
455 290
2 2 3 0 0 0 0 6 3 0 0 3
607 251
642 251
642 276
2 1 5 0 0 4224 0 4 6 0 0 2
534 251
571 251
0
0
25 0 2
0
0
0
0 0 0
0
0 0 0
10000 0 1 10000
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
2689934 1210432 100 100 0 0
0 0 0 0
0 71 161 141
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 0.1
0
396240 8550464 100 100 0 0
77 66 917 396
960 71 1920 560
77 66
917 66
917 66
917 396
0 0
0 0.005 1.2 -1.2 0.005 0.005
12401 0
4 0.001 0.5
2
463 265
0 4 0 0 2	0 4 0 0
621 251
0 3 0 0 1	0 6 0 0
462278 4356672 100 100 0 0
77 66 917 396
958 561 1919 1050
77 66
917 66
917 66
917 330
0 0
1 10000 1.2 0.24 9999 9999
12385 0
4 1000 2000
2
463 271
0 4 0 0 2	0 4 0 0
627 251
0 3 0 0 1	0 6 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
